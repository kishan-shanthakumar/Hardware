module ras
#(parameter ras_size = 8)
(
    input logic clk, rst,
    input logic [63:0] idata,
    output logic [63:0] odata,
    input logic push, pop
);

endmodule