module top(input logic clk, rst,
            output logic trap);

logic [4:0] pipeline_valid;
logic illegal_instr;

endmodule