module wallace_tree_addition #(
    parameter N=32,
    parameter n_products = N*N
) (
    input logic [2*N-1:0] inps [n_products-1:0],
    output logic [2*N-1:0] out
);
genvar i;
generate
    
endgenerate

endmodule