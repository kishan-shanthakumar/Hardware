module stage2(input logic [31:0] instr,
            output [4:0] r1_addr, r2_addr, r3_addr, w1_addr,
            output [3:0] reg_control,
            output [20:0] imm,
            output [1:0] eu_type,
            input clk, rst);

endmodule