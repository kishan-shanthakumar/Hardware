module stage2(input logic [31:0] instr,
            output [4:0] r1_addr, r2_addr, w1_addr,
            // output eu_type,
            input clk, rst);
endmodule