module barrel_shifter(input [63:0] logic op1,
                    input [5:0] logic op2,
                    input logic dir, //1 is left 0 is right
                    output [63:0] logic result);

always_comb
begin

end

endmodule