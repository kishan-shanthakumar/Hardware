module int_div #(parameter N = 32) (
    input logic [N-1:0] a,b,
	output logic [N-1:0] rem,
	output logic [N-1:0] quo
);

endmodule