module stage3();

jumpbranch u1();
base u2();
muldiv u3();

endmodule